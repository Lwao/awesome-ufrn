library verilog;
use verilog.vl_types.all;
entity reg_mult_vlg_vec_tst is
end reg_mult_vlg_vec_tst;
