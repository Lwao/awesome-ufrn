library verilog;
use verilog.vl_types.all;
entity adder_4B_vlg_vec_tst is
end adder_4B_vlg_vec_tst;
