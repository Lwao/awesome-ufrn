library verilog;
use verilog.vl_types.all;
entity parkOmeter_vlg_vec_tst is
end parkOmeter_vlg_vec_tst;
